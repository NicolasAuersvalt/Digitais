	--------------------------------------------------------------------------------
-- Project :
-- File    :
-- Autor   :
-- Date    :
--
--------------------------------------------------------------------------------
-- Description :
--
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Conv_bin_gray IS
  PORT (
  ------------------------------------------------------------------------------
	BIN_IN	: IN std_logic_vector(3 downto 0);
  ------------------------------------------------------------------------------
	GRAY_OUT_VHDL	: OUT std_logic_vector(3 downto 0)
    );
END Conv_bin_gray;

--------------------------------------------------------------------------------
--Complete your VHDL description below
--------------------------------------------------------------------------------

ARCHITECTURE TypeArchitecture OF Conv_bin_gray IS

BEGIN

 ------------------------------------------------------------------------------
	GRAY_OUT_VHDL(3) <=  BIN_IN(3);
	GRAY_OUT_VHDL(2) <= BIN_IN(3) XOR BIN_IN(2);
	GRAY_OUT_VHDL(1) <= BIN_IN(2) XOR BIN_IN(1);
	GRAY_OUT_VHDL(0) <= BIN_IN(1) XOR BIN_IN(0);
 ------------------------------------------------------------------------------	

END TypeArchitecture;
