--------------------------------------------------------------------------------
-- Project :
-- File    :
-- Autor   :
-- Date    :
--
--------------------------------------------------------------------------------
-- Description :
--
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ex_01_a IS
  PORT (
  ------------------------------------------------------------------------------
  --Insert input ports below
    S,R      : IN  std_logic;                    
  ------------------------------------------------------------------------------
  --Insert output ports below
    Q,QN        : OUT std_logic                

    );
END ex_01_a;

--------------------------------------------------------------------------------
--Complete your VHDL description below
--------------------------------------------------------------------------------

ARCHITECTURE TypeArchitecture OF ex_01_a IS
SIGNAL qstate : std_logic;

BEGIN
  PROCESS(S,R)
  BEGIN
    IF (S = '0' AND R = '1') THEN
      qstate <= '1';
    ELSIF (S = '1' AND R = '0') THEN
      qstate <= '0';
    END IF;
  END PROCESS;

  Q <= qstate;
  QN <= NOT qstate;

END TypeArchitecture;
