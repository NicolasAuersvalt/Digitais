LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Aula_03_ex_01 IS
  PORT (
    cnt_i : IN  std_logic_vector(3 downto 0);       -- entrada
    c_7s  : OUT std_logic_vector(6 downto 0)       -- sa�da display
    
  );
END Aula_03_ex_01;

ARCHITECTURE TypeArchitecture OF Aula_03_ex_01 IS
BEGIN

  -- sele��o correta: usa cnt_i, n�o o nome da entidade
  with cnt_i select
    c_7s <= "1111110" when "0000",  -- 0
            "0110000" when "0001",  -- 1
            "1101101" when "0010",  -- 2
            "1111001" when "0011",  -- 3
            "0110011" when "0100",  -- 4
            "1011011" when "0101",  -- 5
            "1011111" when "0110",  -- 6
            "1110000" when "0111",  -- 7
            "1111111" when "1000",  -- 8
            "1110011" when "1001",  -- 9
            "1110111" when "1010",  -- A
            "0011111" when "1011",  -- b
            "1001110" when "1100",  -- C
            "0111101" when "1101",  -- d
            "1011111" when "1110",  -- E
            "1100111" when "1111",  -- F
            "0000000" when others;  -- default (opcional)
            
END TypeArchitecture;
