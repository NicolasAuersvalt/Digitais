--------------------------------------------------------------------------------
-- Project :
-- File    :
-- Autor   :
-- Date    :
--
--------------------------------------------------------------------------------
-- Description :
--
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Aula_02_ex_01 IS
  PORT (
  ------------------------------------------------------------------------------
  --Insert input ports below
    X      : IN  std_logic;                    -- input bit example
    Y      : IN  std_logic;                    -- input bit example
  ------------------------------------------------------------------------------
  --Insert output ports below
    A1        : OUT std_logic;                    -- output bit example
    A2        : OUT std_logic;                    -- output bit example
    B1        : OUT std_logic;                    -- output bit example
    B2        : OUT std_logic                    -- output bit example


    );
END Aula_02_ex_01;

--------------------------------------------------------------------------------
--Complete your VHDL description below
--------------------------------------------------------------------------------

ARCHITECTURE TypeArchitecture OF Aula_02_ex_01 IS

BEGIN
	A1 <= NOT (X OR Y);
	A2 <= (NOT X) AND (NOT Y);
	B1 <= NOT (X AND Y);
	B2 <= (NOT X) OR (NOT Y);
	

END TypeArchitecture;
